module float_point_classify
#(
	parameter FLOAT_POINT_NUMBER_PRECISION = "";
)
(

);



endmodule //float_point_classify
