`include "parameters.h"

module inst_decoder
(
	input [(`INSTS_FETCH_WIDTH_IN_BITS) - 1 : 0]	inst_from_ifetcher_in

);


endmodule
