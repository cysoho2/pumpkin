`ifndef SIMULATION
    `define SIMULATION
    `timescale 100ps/100ps
    `define FULL_CYCLE_DELAY 80
    `define HALF_CYCLE_DELAY 40
    `define MEM_IMAGE_DIR "/Users/pobu/Codes/pumpkin/verify/unit_test/mem_image"
    `define DUMP_FILENAME "sim_waves.fst"
`else
`endif
