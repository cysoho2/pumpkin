`include "sim_config.vh"

`ifndef PARAMETERS
    `define PARAMETERS
    `define BYTE_LEN_IN_BITS                                8
`endif

